/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Paweł Zięba  
 *
 * Description:
 * Package with text configuration.
 */

package text_cfg_pkg;

localparam TEXT_COLOR = 12'h0_0_0;
localparam FONT_RECT_WIDTH = 128;
localparam FONT_RECT_HEIGHT = 256;
localparam CHAR_NUMBER = 256;
localparam CHAR_BIT_LENGTH = 8;
localparam HOR_CHAR_NUMBER = 16;

endpackage
