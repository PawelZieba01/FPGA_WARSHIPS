/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Pawel Zieba
 *
 * Description:
 * Package with confi parameters for background service.
 */

package bg_cfg_pkg;

localparam BORDER_WIDTH = 3;
localparam BACKGROUND_COLOR = 12'hA_A_A;

endpackage
